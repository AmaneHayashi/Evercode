LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY extr_st IS --������״̬����
	PORT(
		clk:           IN STD_LOGIC;
		ISxns:         IN STD_LOGIC; --ʤ��
		ISfail:        IN STD_LOGIC; --ʧ��
		
		statecode:     OUT STD_LOGIC_VECTOR(1 DOWNTO 0) --״̬��
		);
END extr_st;

ARCHITECTURE aextr_st OF extr_st IS 
	
	SIGNAL tempstate:  STD_LOGIC_VECTOR(1 DOWNTO 0);
	
BEGIN 

p1:PROCESS(clk, ISxns, ISfail)
BEGIN 
    IF clk'EVENT AND clk='1' THEN
		IF ISxns ='1' AND ISfail = '0' THEN --ʤ��״̬
			tempstate <="01";
		ELSIF ISfail = '1' AND ISxns = '0' THEN --ʧ��״̬
			tempstate <="10";
		END IF ;
	END IF;
END PROCESS;
	
    statecode<=tempstate;

END aextr_st;
	